module VGA(HS, VS, R, G, B, clk)
{
    output HS,
    output VS,
    output R,
    output G,
    output B,
    input clk
}



endmodule
