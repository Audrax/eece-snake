module LFSR
(
    output bit
);

dff_en dff1
(
    
);

dff_en dff1
(
    
);

dff_en dff1
(
    
);

dff_en dff1
(
    
);

dff_en dff1
(
    
);

dff_en dff1
(
    
);

dff_en dff1
(
    
);

dff_en dff1
(
    
);

dff_en dff1
(
    
);

dff_en dff1
(
    
);

dff_en dff1
(
    
);

dff_en dff1
(
    
);

dff_en dff1
(
    
);

dff_en dff1
(
    
);

dff_en dff1
(
    
);

dff_en dff1
(
    
);
