module collisionDetect
(
    input [19:0] headX, headY, bodyX, bodyY,
    input walls,
    output gameOver
);



endmodule